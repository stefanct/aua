-- ROM file, generated

library ieee;
use ieee.std_logic_1164.all;

entity rom is
port (
		clk : in std_logic;
		address : in std_logic_vector(15 downto 0);
		q : out std_logic_vector(15 downto 0)
);
end rom;

architecture rtl of rom is

signal data : std_logic_vector(15 downto 0);

begin

q <= data;

process(address) begin

	case address is
		when "1000000000000000" => data <= "0110011111100011";	-- addi $3 0x3f
		when "1000000000000010" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000000100" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000000110" => data <= "1100000001000011";	-- lsli $3 2
		when "1000000000001000" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000001010" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000001100" => data <= "0110000001100011";	-- addi $3 3
		when "1000000000001110" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000010000" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000010010" => data <= "1100000100000011";	-- lsli $3 8
		when "1000000000010100" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000010110" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000011000" => data <= "0110001000000011";	-- addi $3 0x10
		when "1000000000011010" => data <= "0110000011000100";	-- addi $4 0x6
		when "1000000000011100" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000011110" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000100000" => data <= "1100000010000100";	-- lsli $4 4
		when "1000000000100010" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000100100" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000100110" => data <= "0110000011000100";	-- addi $4 0x6
		when "1000000000101000" => data <= "1111110010000011";	-- stb $3 $4
		when "1000000000101010" => data <= "0110000010000100";	-- addi $4 0x4
		when "1000000000101100" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000101110" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000110000" => data <= "1100000010000100";	-- lsli $4 4
		when "1000000000110010" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000110100" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000110110" => data <= "0110000111100100";	-- addi $4 0xf
		when "1000000000111000" => data <= "0110000000100011";	-- addi $3 1
		when "1000000000111010" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000111100" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000000111110" => data <= "1111110010000011";	-- stb $3 $4
		when "1000000001000000" => data <= "0110000010100100";	-- addi $4 0x5
		when "1000000001000010" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001000100" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001000110" => data <= "1100000010000100";	-- lsli $4 4
		when "1000000001001000" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001001010" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001001100" => data <= "0110000101100100";	-- addi $4 0xb
		when "1000000001001110" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001010000" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001010010" => data <= "0110000000100011";	-- addi $3 1
		when "1000000001010100" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001010110" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001011000" => data <= "1111110010000011";	-- stb $3 $4
		when "1000000001011010" => data <= "0110000011000100";	-- addi $4 0x06
		when "1000000001011100" => data <= "0110000000100011";	-- addi $3 1
		when "1000000001011110" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001100000" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001100010" => data <= "1111110010000011";	-- stb $3 $4
		when "1000000001100100" => data <= "1100101000100100";	-- scb $4 17
		when "1000000001100110" => data <= "1100101001100010";	-- scb $2 19
		when "1000000001101000" => data <= "1100100001000110";	-- scb $6 2
		when "1000000001101010" => data <= "1100100011100001";	-- scb $1 7
		when "1000000001101100" => data <= "0000000000000000";	-- ldi $0 0
		when "1000000001101110" => data <= "0100000000000000";	-- brezi $0 loop
		when others => data <= "0000000000000000";
	end case;
end process;

end rtl;
