ram_inst : ram PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		rdaddress_a	 => rdaddress_a_sig,
		rdaddress_b	 => rdaddress_b_sig,
		wraddress	 => wraddress_sig,
		wren	 => wren_sig,
		qa	 => qa_sig,
		qb	 => qb_sig
	);
