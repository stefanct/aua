-- Program test/boot.asm, generated ROM file

library ieee;
use ieee.std_logic_1164.all;

entity rom is
port (
		clk : in std_logic;
		address : in std_logic_vector(15 downto 0);
		q : out std_logic_vector(15 downto 0)
);
end rom;

architecture rtl of rom is

signal data : std_logic_vector(15 downto 0);

begin

q <= data;

process(address) begin

	case address is
		when "1000000000000000" => data <= "0000111111111110";	-- 0x8000: ldih $fp, STACK_TOP (ldiw $fp, STACK_TOP)
		when "1000000000000010" => data <= "1100000100011110";	-- 0x8002: lsli $fp, 8 (ldiw $fp, STACK_TOP)
		when "1000000000000100" => data <= "0001111111011110";	-- 0x8004: ldil $fp, STACK_TOP (ldiw $fp, STACK_TOP)
		when "1000000000000110" => data <= "0000111111111101";	-- 0x8006: ldih $sp, STACK_TOP (ldiw $sp, STACK_TOP)
		when "1000000000001000" => data <= "1100000100011101";	-- 0x8008: lsli $sp, 8 (ldiw $sp, STACK_TOP)
		when "1000000000001010" => data <= "0001111111011101";	-- 0x800a: ldil $sp, STACK_TOP (ldiw $sp, STACK_TOP)
		when "1000000000001100" => data <= "0001111111110000";	-- 0x800c: ldih $16, SC_DIGITS (ldiw $16, SC_DIGITS)
		when "1000000000001110" => data <= "1100000100010000";	-- 0x800e: lsli $16, 8 (ldiw $16, SC_DIGITS)
		when "1000000000010000" => data <= "0000001000010000";	-- 0x8010: ldil $16, SC_DIGITS (ldiw $16, SC_DIGITS)
		when "1000000000010010" => data <= "0000000000001010";	-- 0x8012: ldih $10, 0 (ldiw $10, 0)
		when "1000000000010100" => data <= "1100000100001010";	-- 0x8014: lsli $10, 8 (ldiw $10, 0)
		when "1000000000010110" => data <= "0000000000001010";	-- 0x8016: ldil $10, 0 (ldiw $10, 0)
		when "1000000000011000" => data <= "0000000000001011";	-- 0x8018: ldih $11, 1 (ldiw $11, 1)
		when "1000000000011010" => data <= "1100000100001011";	-- 0x801a: lsli $11, 8 (ldiw $11, 1)
		when "1000000000011100" => data <= "0000000000101011";	-- 0x801c: ldil $11, 1 (ldiw $11, 1)
		when "1000000000011110" => data <= "0001000000000010";	-- 0x801e: ldih $2, uart_read (ldiw $2, uart_read)
		when "1000000000100000" => data <= "1100000100000010";	-- 0x8020: lsli $2, 8 (ldiw $2, uart_read)
		when "1000000000100010" => data <= "0000101101000010";	-- 0x8022: ldil $2, uart_read (ldiw $2, uart_read)
		when "1000000000100100" => data <= "1111101110111111";	-- 0x8024: st $ra, $sp (call $2)
		when "1000000000100110" => data <= "0110111111011101";	-- 0x8026: addi $sp, -2 (call $2)
		when "1000000000101000" => data <= "0011010001000000";	-- 0x8028: jmpl $2 (call $2)
		when "1000000000101010" => data <= "0110000001011101";	-- 0x802a: addi $sp, 2 (call $2)
		when "1000000000101100" => data <= "1111001110111111";	-- 0x802c: ld $ra, $sp (call $2)
		when "1000000000101110" => data <= "0001111111100101";	-- 0x802e: ldih $5, SC_DIGITS (ldiw $5, SC_DIGITS)
		when "1000000000110000" => data <= "1100000100000101";	-- 0x8030: lsli $5, 8 (ldiw $5, SC_DIGITS)
		when "1000000000110010" => data <= "0000001000000101";	-- 0x8032: ldil $5, SC_DIGITS (ldiw $5, SC_DIGITS)
		when "1000000000110100" => data <= "0110000000100101";	-- 0x8034: addi $5, 1
		when "1000000000110110" => data <= "0000000000000110";	-- 0x8036: ldih $6, 1 (ldiw $6, 1)
		when "1000000000111000" => data <= "1100000100000110";	-- 0x8038: lsli $6, 8 (ldiw $6, 1)
		when "1000000000111010" => data <= "0000000000100110";	-- 0x803a: ldil $6, 1 (ldiw $6, 1)
		when "1000000000111100" => data <= "1111100010100110";	-- 0x803c: st $6, $5
		when "1000000000111110" => data <= "1111000101001011";	-- 0x803e: ld $11, $10
		when "1000000001000000" => data <= "1111101000001011";	-- 0x8040: st $11, $16
		when "1000000001000010" => data <= "1111101110111111";	-- 0x8042: st $ra, $sp (call $2)
		when "1000000001000100" => data <= "0110111111011101";	-- 0x8044: addi $sp, -2 (call $2)
		when "1000000001000110" => data <= "0011010001000000";	-- 0x8046: jmpl $2 (call $2)
		when "1000000001001000" => data <= "0110000001011101";	-- 0x8048: addi $sp, 2 (call $2)
		when "1000000001001010" => data <= "1111001110111111";	-- 0x804a: ld $ra, $sp (call $2)
		when "1000000001001100" => data <= "0110000000100101";	-- 0x804c: addi $5, 1
		when "1000000001001110" => data <= "0000000000000110";	-- 0x804e: ldih $6, 2 (ldiw $6, 2)
		when "1000000001010000" => data <= "1100000100000110";	-- 0x8050: lsli $6, 8 (ldiw $6, 2)
		when "1000000001010010" => data <= "0000000001000110";	-- 0x8052: ldil $6, 2 (ldiw $6, 2)
		when "1000000001010100" => data <= "1111100010100110";	-- 0x8054: st $6, $5
		when "1000000001010110" => data <= "0000000000000000";	-- 0x8056: ldi $0, 0 (nop)
		when "1000000001011000" => data <= "0011101111100000";	-- 0x8058: brez $0, $31 (ret)
		when "1000000001011010" => data <= "0001111111110100";	-- 0x805a: ldih $20, SC_DIGITS (ldiw $20, SC_DIGITS)
		when "1000000001011100" => data <= "1100000100010100";	-- 0x805c: lsli $20, 8 (ldiw $20, SC_DIGITS)
		when "1000000001011110" => data <= "0000001000010100";	-- 0x805e: ldil $20, SC_DIGITS (ldiw $20, SC_DIGITS)
		when "1000000001100000" => data <= "0000000000010101";	-- 0x8060: ldih $21, 0xf (ldiw $21, 0xf)
		when "1000000001100010" => data <= "1100000100010101";	-- 0x8062: lsli $21, 8 (ldiw $21, 0xf)
		when "1000000001100100" => data <= "0000000111110101";	-- 0x8064: ldil $21, 0xf (ldiw $21, 0xf)
		when "1000000001100110" => data <= "1111101010010101";	-- 0x8066: st $21, $20
		when "1000000001101000" => data <= "1111101110100001";	-- 0x8068: st $1, $sp (push $1)
		when "1000000001101010" => data <= "0110111111011101";	-- 0x806a: addi $sp, -2 (push $1)
		when "1000000001101100" => data <= "1111101110100010";	-- 0x806c: st $2, $sp (push $2)
		when "1000000001101110" => data <= "0110111111011101";	-- 0x806e: addi $sp, -2 (push $2)
		when "1000000001110000" => data <= "1111101110100011";	-- 0x8070: st $3, $sp (push $3)
		when "1000000001110010" => data <= "0110111111011101";	-- 0x8072: addi $sp, -2 (push $3)
		when "1000000001110100" => data <= "1111101110100100";	-- 0x8074: st $4, $sp (push $4)
		when "1000000001110110" => data <= "0110111111011101";	-- 0x8076: addi $sp, -2 (push $4)
		when "1000000001111000" => data <= "1111101110101010";	-- 0x8078: st $10, $sp (push $10)
		when "1000000001111010" => data <= "0110111111011101";	-- 0x807a: addi $sp, -2 (push $10)
		when "1000000001111100" => data <= "1111101110101011";	-- 0x807c: st $11, $sp (push $11)
		when "1000000001111110" => data <= "0110111111011101";	-- 0x807e: addi $sp, -2 (push $11)
		when "1000000010000000" => data <= "0001111111100001";	-- 0x8080: ldih $1, SC_UART_STATUS (ldiw $1, SC_UART_STATUS)
		when "1000000010000010" => data <= "1100000100000001";	-- 0x8082: lsli $1, 8 (ldiw $1, SC_UART_STATUS)
		when "1000000010000100" => data <= "0000010000000001";	-- 0x8084: ldil $1, SC_UART_STATUS (ldiw $1, SC_UART_STATUS)
		when "1000000010000110" => data <= "0001111111100100";	-- 0x8086: ldih $4, SC_UART_DATA (ldiw $4, SC_UART_DATA)
		when "1000000010001000" => data <= "1100000100000100";	-- 0x8088: lsli $4, 8 (ldiw $4, SC_UART_DATA)
		when "1000000010001010" => data <= "0000010000100100";	-- 0x808a: ldil $4, SC_UART_DATA (ldiw $4, SC_UART_DATA)
		when "1000000010001100" => data <= "0000000000100011";	-- 0x808c: ldi $3, 1
		when "1000000010001110" => data <= "1111000000100010";	-- 0x808e: ld $2, $1
		when "1000000010010000" => data <= "1010010001000011";	-- 0x8090: and $3, $2
		when "1000000010010010" => data <= "0100111110100011";	-- 0x8092: brezi $3, loop_read
		when "1000000010010100" => data <= "1111000010000010";	-- 0x8094: ld $2, $4
		when "1000000010010110" => data <= "1111100101000010";	-- 0x8096: st $2, $10
		when "1000000010011000" => data <= "0001111111100101";	-- 0x8098: ldih $5, SC_DIGITS (ldiw $5, SC_DIGITS)
		when "1000000010011010" => data <= "1100000100000101";	-- 0x809a: lsli $5, 8 (ldiw $5, SC_DIGITS)
		when "1000000010011100" => data <= "0000001000000101";	-- 0x809c: ldil $5, SC_DIGITS (ldiw $5, SC_DIGITS)
		when "1000000010011110" => data <= "1111100010100010";	-- 0x809e: st $2, $5
		when "1000000010100000" => data <= "0110000001001010";	-- 0x80a0: addi $10, 2
		when "1000000010100010" => data <= "0110111111101011";	-- 0x80a2: addi $11, -1
		when "1000000010100100" => data <= "0101111010001011";	-- 0x80a4: brnezi $11, loop_read
		when "1000000010100110" => data <= "0110000001011101";	-- 0x80a6: addi $sp, 2 (pop $11)
		when "1000000010101000" => data <= "1111001110101011";	-- 0x80a8: ld $11, $sp (pop $11)
		when "1000000010101010" => data <= "0110000001011101";	-- 0x80aa: addi $sp, 2 (pop $10)
		when "1000000010101100" => data <= "1111001110101010";	-- 0x80ac: ld $10, $sp (pop $10)
		when "1000000010101110" => data <= "0110000001011101";	-- 0x80ae: addi $sp, 2 (pop $4)
		when "1000000010110000" => data <= "1111001110100100";	-- 0x80b0: ld $4, $sp (pop $4)
		when "1000000010110010" => data <= "0110000001011101";	-- 0x80b2: addi $sp, 2 (pop $3)
		when "1000000010110100" => data <= "1111001110100011";	-- 0x80b4: ld $3, $sp (pop $3)
		when "1000000010110110" => data <= "0110000001011101";	-- 0x80b6: addi $sp, 2 (pop $2)
		when "1000000010111000" => data <= "1111001110100010";	-- 0x80b8: ld $2, $sp (pop $2)
		when "1000000010111010" => data <= "0110000001011101";	-- 0x80ba: addi $sp, 2 (pop $1)
		when "1000000010111100" => data <= "1111001110100001";	-- 0x80bc: ld $1, $sp (pop $1)
		when "1000000010111110" => data <= "0011101111100000";	-- 0x80be: brez $0, $31 (ret)
		when "1000000110000000" => data <= "0000000001000000";
		when "1000000110000010" => data <= "0000000001111001";
		when "1000000110000100" => data <= "0000000000100100";
		when "1000000110000110" => data <= "0000000000110000";
		when "1000000110001000" => data <= "0000000000011001";
		when "1000000110001010" => data <= "0000000000010010";
		when "1000000110001100" => data <= "0000000000000010";
		when "1000000110001110" => data <= "0000000001111000";
		when "1000000110010000" => data <= "0000000000000000";
		when "1000000110010010" => data <= "0000000000010000";
		when others => data <= "0000000000000000";
	end case;
end process;

end rtl;
